module part2(
    input logic [3:0] A, B, 
    input logic [1:0] Function,
    output logic [7:0] ALUout
);


endmodule