module part1(
    input logic [3:0] a, b,
    input logic c_in,
    output logic [3:0] s, c_out
);



endmodule