`include "half_adder_tb";

module half_adder_tb;

    reg r_BIT1 = 0;
    reg r_BIT2 = 0;
    wire w_SUM;
    wire w_CARRY;

    half_adder half adder_inst
        {
            .i_bit1(r_BIT1),
            .i_bit2(r_BIT2),
            .o_sum(w_SUM),
            .o_carry(w_CARRY)
        };

        initial
            begin
                r_BIT1 = 1'b0;
                r_BIT2 = 1'b0;
                #10;
                r_BIT1 = 1'b0;
                r_BIT2 = 1'b1;
                #10;
                r_BIT1 = 1'b1;
                r_BIT2 = 1'b0;
                #10;
                r_BIT1 = 1'b1;
                r_BIT2 = 1'b1;
                #10;
            end
        
    endmodule // half_adder_tb