module part2
#(parameter CLOCK_FREQUENCY=500)(
    input logic ClockIn, Reset,
    input logic [1:0] Speed,
    output logic [3:0] CounterValue
);

endmodule