`include "Full_Adder.v"

module carry_lookahead_adder_4_bit
    (
        input [3:0]     i_add1,
        input [3:0]     i_add2,
        output [4:0]    o_result
    );

    wire [4:0]      w_C;
    wire [3:0]      w_G, w_P, w_SUM;

    full_adder full_adder_bit_0
        (
            .i_bit1(i_add1[0]),
            .i_bit2(i_add2[0]),
            .i_carry(w_C[0]),    
            .o_sum(w_SUM[0]),
            .o_carry()   
        );

    full_adder full_adder_bit_1
        (
            .i_bit1(i_add1[1]),
            .i_bit2(i_add2[1]),
            .i_carry(w_C[1]),    
            .o_sum(w_SUM[1]),
            .o_carry()   
        );

    full_adder full_adder_bit_2
        (
            .i_bit1(i_add1[2]),
            .i_bit2(i_add2[2]),
            .i_carry(w_C[2]),    
            .o_sum(w_SUM[2]),
            .o_carry()   
        );

    full_adder full_adder_bit_3
        (
            .i_bit1(i_add1[3]),
            .i_bit2(i_add2[3]),
            .i_carry(w_C[3]),    
            .o_sum(w_SUM[3]),
            .o_carry()   
        );

    // Create the Generate (G) Terms: G_i = A_i * B_i
    assign w_G[0] = i_add1[0] & i_add2[0];
    assign w_G[1] = i_add1[1] & i_add2[1];
    assign w_G[2] = i_add1[2] & i_add2[2];
    assign w_G[3] = i_add1[3] & i_add2[3];

    // Create the Propagate Terms: P_i = A_i + B_i
    assign w_P[0] = i_add1[0] & i_add2[0];
    assign w_P[1] = i_add1[1] & i_add2[1];
    assign w_P[2] = i_add1[2] & i_add2[2];
    assign w_P[3] = i_add1[3] & i_add2[3];
    
    // Creat the Carry Terms:
    assign w_C[0] = 1'b0 // no carry input
    assign w_C[1] = w_G[1] | (w_P[1] & w_C[1]);
    assign w_C[2] = w_G[2] | (w_P[2] & w_C[2]);
    assign w_C[3] = w_G[3] | (w_P[3] & w_C[3]);
    assign w_C[4] = w_G[4] | (w_P[4] & w_C[4]);

    assign i_result = {w_C[4], w_SUM}; // Verilog Concatentation

endmodule // carry_lookahead_adder_4_bit