module part3(
    input logic Clock, Reset_b,
    input logic [3:0] Data,
    input logic [2:0] Function,
    output logic [7:0] ALU_reg_out
);

endmodule