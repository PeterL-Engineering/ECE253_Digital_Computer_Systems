module part3
#(parameter CLOCK_FREQUENCY=500)(
    input logic ClockIn, Reset, Start,
    input logic [2:0] Letter,
    output logic DotDashOut, NewBitOu
);

endmodule