module part1(
    input logic clock, reset, ParallelLoadn, RotateRight, ASRight,
    input logic [3:0] Data_IN,
    output logic [3:0] Q
);

endmodule